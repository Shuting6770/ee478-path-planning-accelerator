`define FSB_LEGACY
